`ifndef BRAM_A_SEQ_LIB_SV
`define BRAM_A_SEQ_LIB_SV

`include "bram_a_basic_seq.sv"

`endif // BRAM_A_SEQ_LIB_SV
