`ifndef AXI_LITE_SEQ_LIB_SV
`define AXI_LITE_SEQ_LIB_SV

`include "axi_lite_basic_seq.sv"
`include "axi_lite_write_start_register_value_seq.sv"
`include "axi_lite_read_ready_register_seq.sv"



`endif // AXI_LITE_SEQ_LIB_SV
